package shared_pkg;
    int error_count;
    int all_error_count;
    int correct_count;
    int all_correct_count;
    bit test_finished;
    event input_driven;
endpackage